library ieee;
use ieee.std_logic_1164.all;

entity zeroextend is
	port(input: in std_logic_vector(8 downto 0);
		  output: out std_logic_vector(15 downto 0));
end entity;

architecture zeroarch of zeroextend is

begin
	extend_7: process(input)
	
	
	begin
		output(8 downto 0) <= input;
		output(15 downto 9) <= "0000000";

	end process;
		
		
end zeroarch;