-- THIS IS THE CODE FOR THE ARF AND RRF
library ieee;
use ieee.std_logic_1164.all;

entity ARF is
	port(opr1, opr2,opr3: in std_logic_vector(2 downto 0);
	clk , rst  : in std_logic;
	
	)